`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/30/2024 03:40:48 PM
// Design Name: 
// Module Name: InstructionsMemory
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module InstructionsMemory(
    input [31:0] Address,
    output reg [31:0] Instructions
    );
    
always @(*) begin
    case(Address)
//*********************************A PROGRAM CHECKS HAZARDS&JAL&JALR INSTRUCTIONS*********************************
//    32'h00000000: Instructions = 32'b00000000000100000000000010010011; // 	  addi x1, x0, 1 //0
//    32'h00000004: Instructions = 32'b00000000000100000000000100110011; // 	  add x2, x0, x1 //4 
//    32'h00000008: Instructions = 32'b00000000001000000010000000100011; // 	  sw  x2 ,0(x0)  // 8
//    32'h0000000c: Instructions = 32'b00000000000000000010000110000011; // 	  lw  x3 ,0(x0)  //12
//    32'h00000010: Instructions = 32'b00000000000100000000001000010011; // 	  addi x4, x0, 1 // 16
//    32'h00000014: Instructions = 32'b00000000001000100000100001100011; // 	  beq  x4, x2, check_beq //20
//    32'h00000018: Instructions = 32'b00000000000100000000001100010011; //       addi x6, x0, 1 //24
//    32'h0000001c: Instructions = 32'b00000000000100000000001100010011; //       addi x6, x0, 1 //28
//    32'h00000020: Instructions = 32'b00000000000100000000001100010011; //       addi x6, x0, 1 //32
//    32'h00000024: Instructions = 32'b00000000000100000000001010010011; // 	  check_beq:	addi x5, x0, 1 //36
//    32'h00000028: Instructions = 32'b00000000000000000010010010000011; // 	  lw   x9, 0(x0) //40 
//    32'h0000002c: Instructions = 32'b00000000011101001000010000110011; //       add  x8, x9, x7 //44
//    32'h00000030: Instructions = 32'b00000000100000000000011001101111; //       jal  x12, check_jal //48
//    32'h00000034: Instructions = 32'b00000000000100000000001100010011; //       addi x6, x0, 1 //52
//    32'h00000038: Instructions = 32'b00000000001000000000001100010011; //       check_jal:	addi x6, x0, 2 //56
//    32'h0000003c: Instructions = 32'b00000100000000000000001110010011; //       addi x7, x0, 0x40 //60
//    32'h00000040: Instructions = 32'b00000000110000111000010111100111; //       jalr x11, x7, 0xc //64
//    32'h00000044: Instructions = 32'b00000000000100000000010100010011; //       addi x10, x0, 1 //68
//    32'h00000048: Instructions = 32'b00000000001000000000010100010011; //       addi x10, x0, 2 //72
//    32'h0000004c: Instructions = 32'b00000000001100000000010100010011; //       addi x10, x0, 3 //76
    
//*********************************A PROGRAM CHECKS LOAD&STORE INSTRUCTIONS*********************************  
//    32'h00000000: Instructions = 32'b11111111111100000000000010010011; // 	addi x1, x0, 0xfff
//    32'h00000004: Instructions = 32'b00000000000100000010000000100011; // 	sw   x1, 0(x0)
//    32'h00000008: Instructions = 32'b00000000000000000010000100000011; // 	lw   x2, 0(x0)
//    32'h0000000c: Instructions = 32'b00000000000000000000000110000011; // 	lb   x3, 0(x0)
//    32'h00000010: Instructions = 32'b00000000000000000001001000000011; // 	lh   x4, 0(x0)
//    32'h00000014: Instructions = 32'b00000000000000000100001010000011; // 	lbu  x5, 0(x0)
//    32'h00000018: Instructions = 32'b00000000000000000101001100000011; //     lhu  x6, 0(x0)
//    32'h0000001c: Instructions = 32'b00000000000100000001001000100011; //     sh   x1, 4(x0)                
//    32'h000000020: Instructions = 32'b00000000000100000000010000100011; //    sb   x1, 8(x0  
             
//*********************************A PROGRAM CHECKS BRANCH INSTRUCTIONS*********************************      
//    32'h00000000: Instructions = 32'b00000000000100000000000010010011; // 	  addi x1, x0, 1
//    32'h00000004: Instructions = 32'b00000000000100000000000100010011; // 	  addi x2, x0, 1
//    32'h00000008: Instructions = 32'b00000000001000000000000110010011; // 	  addi x3, x0, 2
//    32'h0000000c: Instructions = 32'b11111111111100000000111100010011; // 	  addi x30, x0, -1
//    32'h00000010: Instructions = 32'b00000000001100010001010001100011; // 	  bne  x2, x3, check_bne
//    32'h00000014: Instructions = 32'b00000000000100000000001010010011; // 	  addi x5, x0, 1
//    32'h00000018: Instructions = 32'b00000000001000000000001010010011; //     check_bne: addi x5, x0, 2
//    32'h0000001c: Instructions = 32'b00000000001000001000010001100011; //     beq  x1, x2, check_beq
//    32'h00000020: Instructions = 32'b00000000000100000000001000010011; //     addi x4, x0, 1
//    32'h00000024: Instructions = 32'b00000000001000000000001000010011; // 	  check_beq: addi x4, x0, 2
//    32'h00000028: Instructions = 32'b00000000001100010100010001100011; // 	  blt x2, x3, check_blt
//    32'h0000002c: Instructions = 32'b00000000000100000000001100010011; //     addi x6, x0, 1
//    32'h00000030: Instructions = 32'b00000000001000000000001100010011; //     check_blt: addi x6, x0, 2
//    32'h00000034: Instructions = 32'b00000000001000001101010001100011; //     bge  x1, x2, check_bge
//    32'h00000038: Instructions = 32'b00000000000100000000001110010011; //     addi x7, x0, 1
//    32'h0000003c: Instructions = 32'b00000000001000000000001110010011; //     check_bge: addi x7, x0, 2
//    32'h00000040: Instructions = 32'b11111111111100000000111110010011; //     addi x31, x0, -1
//    32'h00000044: Instructions = 32'b00000001111100001111010001100011; //     bgeu x1, x31, check_bgeu
//    32'h00000048: Instructions = 32'b00000000000100000000010000010011; //     addi x8, x0, 1
//    32'h0000004c: Instructions = 32'b00000000001000000000010000010011; //     check_bgeu: addi x8, x0, 2
//    32'h00000050: Instructions = 32'b00000001111000000110010001100011; //     bltu x0, x30, check_bltu
//    32'h00000054: Instructions = 32'b00000000000100000000010010010011; //     addi x9, x0, 1
//    32'h00000058: Instructions = 32'b00000000001000000000010010010011; //     check_bltu: addi x9, x0, 2

//*********************************A PROGRAM CHECKS Itype INSTRUCTIONS********************************* 
//    32'h00000000: Instructions = 32'b00000000001000000000000010010011; // 	  addi x1, x0, 2
//    32'h00000004: Instructions = 32'b00000000001000000000000100010011; // 	  addi x2, x0, 2
//    32'h00000008: Instructions = 32'b00000000000000000001000110110111; // 	  lui  x3, 0x1
//    32'h0000000c: Instructions = 32'b00000000000000000001001000010111; // 	  auipc x4, 0x1
//    32'h00000010: Instructions = 32'b00000000001100001111001010010011; // 	  andi  x5, x1, 3
//    32'h00000014: Instructions = 32'b00000000001100001100001100010011; // 	  xori  x6, x1, 3
//    32'h00000018: Instructions = 32'b00000000001100001110011000010011; //     ori   x12, x1, 3
//    32'h0000001c: Instructions = 32'b00000000001100001010001110010011; //     slti  x7, x1, 3
//    32'h00000020: Instructions = 32'b11111111110100001011010000010011; //     sltiu x8, x1, -3
//    32'h00000024: Instructions = 32'b00000000000100001001010010010011; // 	  slli  x9, x1, 1
//    32'h00000028: Instructions = 32'b00000000000100001101010100010011; // 	  srli  x10, x1, 1
//    32'h0000002c: Instructions = 32'b01000000000100001101010110010011; //     srai  x11, x1, 1

//*********************************A PROGRAM CHECKS Rtype INSTRUCTIONS********************************* 
    32'h00000000: Instructions = 32'b00000000001000000000000010010011; // 	  addi x1, x0, 2
    32'h00000004: Instructions = 32'b00000000000000001000000100110011; // 	  add x2, x1, x0	
    32'h00000008: Instructions = 32'b00000000001000001111000110110011; // 	  and x3, x1, x2
    32'h0000000c: Instructions = 32'b01000000000000001000001000110011; // 	  sub x4, x1, x0
    32'h00000010: Instructions = 32'b00000000001000001001001010110011; //     sll x5, x1, x2
    32'h00000014: Instructions = 32'b00000000010100100010001100110011; //     slt x6, x4, x5
    32'h00000018: Instructions = 32'b11111111110100000000001110010011; //     addi x7, x0, -3
    32'h0000001c: Instructions = 32'b00000000011100001011010000110011; //     sltu x8, x1, x7
    32'h00000020: Instructions = 32'b00000000000100101110010010110011; //     or   x9, x5, x1
    32'h00000024: Instructions = 32'b00000000001000001101010100110011; //     srl  x10, x1, x2
    32'h00000028: Instructions = 32'b01000000001000001101010110110011; //     sra  x11, x1, x2
default: Instructions = 32'dz; 
    
    endcase

end

endmodule
